module or_gate(out, A, B); 

    output [31:0] out;
    input [31:0] A, B; 

    
    or OR0(out[0], A[0], B[0]);
    or OR1(out[1], A[1], B[1]);
    or OR2(out[2], A[2], B[2]);
    or OR3(out[3], A[3], B[3]);
    or OR4(out[4], A[4], B[4]);
    or OR5(out[5], A[5], B[5]);
    or OR6(out[6], A[6], B[6]);
    or OR7(out[7], A[7], B[7]);
    or OR8(out[8], A[8], B[8]);
    or OR9(out[9], A[9], B[9]);
    or OR10(out[10], A[10], B[10]);
    or OR11(out[11], A[11], B[11]);
    or OR12(out[12], A[12], B[12]);
    or OR13(out[13], A[13], B[13]);
    or OR14(out[14], A[14], B[14]);
    or OR15(out[15], A[15], B[15]);
    or OR16(out[16], A[16], B[16]);
    or OR17(out[17], A[17], B[17]);
    or OR18(out[18], A[18], B[18]);
    or OR19(out[19], A[19], B[19]);
    or OR20(out[20], A[20], B[20]);
    or OR21(out[21], A[21], B[21]);
    or OR22(out[22], A[22], B[22]);
    or OR23(out[23], A[23], B[23]);
    or OR24(out[24], A[24], B[24]);
    or OR25(out[25], A[25], B[25]);
    or OR26(out[26], A[26], B[26]);
    or OR27(out[27], A[27], B[27]);
    or OR28(out[28], A[28], B[28]);
    or OR29(out[29], A[29], B[29]);
    or OR30(out[30], A[30], B[30]);
    or OR31(out[31], A[31], B[31]);
endmodule 