module not_bit(result, operand);

    input [31:0] operand;
    output [31:0] result;

    not NOT0(result[0], operand[0]);
    not NOT1(result[1], operand[1]);
    not NOT2(result[2], operand[2]);
    not NOT3(result[3], operand[3]);
    not NOT4(result[4], operand[4]);
    not NOT5(result[5], operand[5]);
    not NOT6(result[6], operand[6]);
    not NOT7(result[7], operand[7]);
    not NOT8(result[8], operand[8]);
    not NOT9(result[9], operand[9]);
    not NOT10(result[10], operand[10]);
    not NOT11(result[11], operand[11]);
    not NOT12(result[12], operand[12]);
    not NOT13(result[13], operand[13]);
    not NOT14(result[14], operand[14]);
    not NOT15(result[15], operand[15]);
    not NOT16(result[16], operand[16]);
    not NOT17(result[17], operand[17]);
    not NOT18(result[18], operand[18]);
    not NOT19(result[19], operand[19]);
    not NOT20(result[20], operand[20]);
    not NOT21(result[21], operand[21]);
    not NOT22(result[22], operand[22]);
    not NOT23(result[23], operand[23]);
    not NOT24(result[24], operand[24]);
    not NOT25(result[25], operand[25]);
    not NOT26(result[26], operand[26]);
    not NOT27(result[27], operand[27]);
    not NOT28(result[28], operand[28]);
    not NOT29(result[29], operand[29]);
    not NOT30(result[30], operand[30]);
    not NOT31(result[31], operand[31]);

endmodule