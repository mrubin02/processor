module bypass_ctrl(select, ir_x, ir_m, ir_w);

    input [31:0] ir_x, ir_m, ir_w;
    output [1:0] select;

    

endmodule