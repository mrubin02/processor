module not_gate(out, A); 
    input [31:0] A; 
    output [31:0] out;

    not NOT0(out[0], A[0]);
    not NOT1(out[1], A[1]);
    not NOT2(out[2], A[2]);
    not NOT3(out[3], A[3]);
    not NOT4(out[4], A[4]);
    not NOT5(out[5], A[5]);
    not NOT6(out[6], A[6]);
    not NOT7(out[7], A[7]);
    not NOT8(out[8], A[8]);
    not NOT9(out[9], A[9]);
    not NOT10(out[10], A[10]);
    not NOT11(out[11], A[11]);
    not NOT12(out[12], A[12]);
    not NOT13(out[13], A[13]);
    not NOT14(out[14], A[14]);
    not NOT15(out[15], A[15]);
    not NOT16(out[16], A[16]);
    not NOT17(out[17], A[17]);
    not NOT18(out[18], A[18]);
    not NOT19(out[19], A[19]);
    not NOT20(out[20], A[20]);
    not NOT21(out[21], A[21]);
    not NOT22(out[22], A[22]);
    not NOT23(out[23], A[23]);
    not NOT24(out[24], A[24]);
    not NOT25(out[25], A[25]);
    not NOT26(out[26], A[26]);
    not NOT27(out[27], A[27]);
    not NOT28(out[28], A[28]);
    not NOT29(out[29], A[29]);
    not NOT30(out[30], A[30]);
    not NOT31(out[31], A[31]);
endmodule 
